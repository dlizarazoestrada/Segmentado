module ex_rurs1(
    input logic clk,
    input logic rst,
    input logic [31:0] ex_rurs1_in = 32'b0, 
    output logic [31:0] ex_rurs1_out
     
);

    always_ff @(posedge clk or negedge rst) begin
        if (rst) begin
            ex_rurs1_out <= 32'b0; 
        end else begin
            ex_rurs1_out <= ex_rurs1_in; 
        end
    end
endmodule